`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:59:07 11/14/2012 
//
//////////////////////////////////////////////////////////////////////////////////
module camera_ctrlr (
	input 			osc_clk_100_bufd,
	input 			clk_50,			// 50Mhz memory clock
	input 			reset,
	// Camera interface
	inout 			CAMA_SDA,
	inout 			CAMA_SCL,
	input 	[7:0] 	CAMA_D_I,
	inout 			CAMA_PCLK_I,
	output 			CAMA_MCLK_O,
	input 			CAMA_LV_I,
	input 			CAMA_FV_I,
	output 			CAMA_RST_O, 	
	output 			CAMA_PWDN_O, 	
	output 			CAMX_VDDEN_O,	
	// Memory interface
	input 			op_begun,
	input			data_ok,
	input 			ctrlr_good,
	output 			mem_wr,
	output 			mem_burst,
	output [15:0] 	mem_data,
	output [22:0] 	mem_addr
	);

wire [15:0] CamAD;

dcm_24_24i dcm_24_24i_inst
(
    .CLK_IN1 		(osc_clk_100_bufd),
    .CLK_24 		(CamClk),
    .CLK_24_inv		(CamClk_180),
    .RESET 			(reset)
);

camera_buffer camera_buffer_inst
(
	// inputs
	.mem_clk 		(clk_50),
	.cam_clk 		(CamAPClk),
	.reset 			(reset),
	.cam_data 		(CAMA_D_I),//(CamAD),
	.cam_fv 		(CAMA_FV_I),
	.cam_lv 		(CAMA_LV_I),
	.op_begun 		(op_begun),
	.data_ok 		(data_ok),
	.ctrlr_good 	(ctrlr_good),
	// outputs
	.mem_wr			(mem_wr),
	.mem_burst		(mem_burst),
	.mem_data		(mem_data),
	.mem_addr		(mem_addr)
);

CamCtl CamCtl_vhdl_inst
(
	.D_O 		(CamAD),				// 15:0 pixel sent to buffer
	.PCLK_O		(CamAPClk),				// buf'd pixel clock (use in fifo)
	.DV_O 		(CamADV),				// pixel data byte select
	.RST_I 		(reset),				// async reset
	.CLK 		(CamClk),				// 24 Mhz controller clock
	.CLK_180 	(CamClk_180),			// 24 Mhz inv controller clock
	.SDA 		(CAMA_SDA),				// inout pin
	.SCL 		(CAMA_SCL),				// inout pin
	.D_I 		(CAMA_D_I),				// 7:0 data from camera (half pixel at a time)
	.PCLK_I 	(int_CAMA_PCLK_I),		// iobuf'd pixel clock generated by camera
	.MCLK_O 	(CAMA_MCLK_O),			// mclk sent to camera (oddr'd in CamCtl)
	.LV_I 		(CAMA_LV_I),			// line valid
	.FV_I 		(CAMA_FV_I),			// frame valid
	.RST_O 		(CAMA_RST_O),			// Reset active LOW
	.PWDN_O 	(CAMA_PWDN_O),			// Power-down active HIGH
	.VDDEN_O 	(CAMX_VDDEN_O)			// common power supply enable (can do power cycle)
);

IOBUF 
#(
 	.DRIVE		(12),
	.IOSTANDARD ("DEFAULT"),
	.SLEW		("SLOW")
)
Inst_IOBUF_CAMA_PCLK 
(
	.O 			(int_CAMA_PCLK_I),  // Buffer output
	.IO 		(CAMA_PCLK_I),   	// Buffer inout port (connect directly to top-level port)
	.I  		(1'b0),     		// Buffer input
	.T 			(1'b1)		      	// 3-state enable input, high=input, low=output 
);

endmodule
